//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_8_x49(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'h00EA1900E5000800F7A0110058000000564A000002000000A9000000B7000000),
.INIT_01(256'h7DAC30009A4623007E391300D3990000B2952900E4DF2B00B9000200A5000000),
.INIT_02(256'hC06E8400A100950037248C001C009D000BCE0000DB000000F48400006E000000),
.INIT_03(256'hF19ECE99A2C0EDA97C8563176591402784806DBE667E5F8E019BC830A92FFA00),
.INIT_04(256'hD0EE6B429A25D56339049F0018A4000041891121BAE2BE00C3008E0053000000),
.INIT_05(256'hB6B35959FE78E578B09D9D00933D0000BE4D233A47268E1BD3008C0041000000),
.INIT_06(256'h278E7F18E9C1C139943ED100311A4E002BE9987B5406375AF33A5D00E7BED300),
.INIT_07(256'h5F377CC8A348F0D98DCD6C451AD9C175EDEEBC8CA031219D5477C76272C37B52),
.INIT_08(256'hFB11E2FB1EFBF3FB0C5BEAFBA3FBFBFBADB1FBFBF9FBFBFB52FBFBFB4CFBFBFB),
.INIT_09(256'h8657CBFB61BDD8FB85C2E8FB2862FBFB496ED2FB1F24D0FB42FBF9FB5EFBFBFB),
.INIT_0A(256'h3B957FFB5AFB6EFBCCDF77FBE7FB66FBF035FBFB20FBFBFB0F7FFBFB95FBFBFB),
.INIT_0B(256'h0A653562593B1652877E98EC9E6ABBDC7F7B96459D85A475FA6033CB52D401FB),
.INIT_0C(256'h2B1590B961DE2E98C2FF64FBE35FFBFBBA72EADA411945FB38FB75FBA8FBFBFB),
.INIT_0D(256'h4D48A2A205831E834B6666FB68C6FBFB45B6D8C1BCDD75E028FB77FBBAFBFBFB),
.INIT_0E(256'hDC7584E3123A3AC26FC52AFBCAE1B5FBD0126380AFFDCCA108C1A6FB1C4528FB),
.INIT_0F(256'hA4CC873358B30B22763697BEE1223A8E161547775BCADA66AF8C3C99893880A9),
.INIT_10(256'h095BAC0045002900165E85005F00000059050000CE0000006F000000FD000000),
.INIT_11(256'hD7AEB5007FF5D400D9476100741900009EE91900EDECFD00B900E400CF000000),
.INIT_12(256'h03FFE000EB0065001CFAC900F1004C001FA100002C00000029A400001F000000),
.INIT_13(256'hECDDC7D8B270F48A16C0E72C4D68D47E97E459A61217EFF444F95052C40FE600),
.INIT_14(256'h51255CF8B31A779C34984F00B7C600005B216C646240C2008B00CA00D3000000),
.INIT_15(256'h4C13863B4A2C495FFB81AB009CDF00005F0EB6A7826FFCC35D002E00E1000000),
.INIT_16(256'h1EDC3ACA584711AE49531B006EA9540058D84656C51DE832BACBD200466F1800),
.INIT_17(256'h2629CAC5D6E057F3577D2138C6D5D86A074AC8272CDDD011C38296468974EA14),
.INIT_18(256'hF2A057FBBEFBD2FBEDA57EFBA4FBFBFBA2FEFBFB35FBFBFB94FBFBFB06FBFBFB),
.INIT_19(256'h2C554EFB840E2FFB22BC9AFB8FE2FBFB6512E2FB161706FB42FB1FFB34FBFBFB),
.INIT_1A(256'hF8041BFB10FB9EFBE70132FB0AFBB7FBE45AFBFBD7FBFBFBD25FFBFBE4FBFBFB),
.INIT_1B(256'h17263C23498B0F71ED3B1CD7B6932F856C1FA25DE9EC140FBF02ABA93FF41DFB),
.INIT_1C(256'hAADEA70348E18C67CF63B4FB4C3DFBFBA0DA979F99BB39FB70FB31FB28FBFBFB),
.INIT_1D(256'hB7E87DC0B1D7B2A4007A50FB6724FBFBA4F54D5C79940738A6FBD5FB1AFBFBFB),
.INIT_1E(256'hE527C131A3BCEA55B2A8E0FB9552AFFBA323BDAD3EE613C9413029FBBD94E3FB),
.INIT_1F(256'hDDD2313E2D1BAC08AC86DAC33D2E2391FCB133DCD7262BEA38796DBD728F11EF),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
	.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
