//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_8_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'h095BAC0045002900165E85005F00000059050000CE0000006F000000FD000000),
.INIT_01(256'hD7AEB5007FF5D400D9476100741900009EE91900EDECFD00B900E400CF000000),
.INIT_02(256'h03FFE000EB0065001CFAC900F1004C001FA100002C00000029A400001F000000),
.INIT_03(256'hECDDC7D8B270F48A16C0E72C4D68D47E97E459A61217EFF444F95052C40FE600),
.INIT_04(256'h51255CF8B31A779C34984F00B7C600005B216C646240C2008B00CA00D3000000),
.INIT_05(256'h4C13863B4A2C495FFB81AB009CDF00005F0EB6A7826FFCC35D002E00E1000000),
.INIT_06(256'h1EDC3ACA584711AE49531B006EA9540058D84656C51DE832BACBD200466F1800),
.INIT_07(256'h2629CAC5D6E057F3577D2138C6D5D86A074AC8272CDDD011C38296468974EA14),
.INIT_08(256'hF2A057FBBEFBD2FBEDA57EFBA4FBFBFBA2FEFBFB35FBFBFB94FBFBFB06FBFBFB),
.INIT_09(256'h2C554EFB840E2FFB22BC9AFB8FE2FBFB6512E2FB161706FB42FB1FFB34FBFBFB),
.INIT_0A(256'hF8041BFB10FB9EFBE70132FB0AFBB7FBE45AFBFBD7FBFBFBD25FFBFBE4FBFBFB),
.INIT_0B(256'h17263C23498B0F71ED3B1CD7B6932F856C1FA25DE9EC140FBF02ABA93FF41DFB),
.INIT_0C(256'hAADEA70348E18C67CF63B4FB4C3DFBFBA0DA979F99BB39FB70FB31FB28FBFBFB),
.INIT_0D(256'hB7E87DC0B1D7B2A4007A50FB6724FBFBA4F54D5C79940738A6FBD5FB1AFBFBFB),
.INIT_0E(256'hE527C131A3BCEA55B2A8E0FB9552AFFBA323BDAD3EE613C9413029FBBD94E3FB),
.INIT_0F(256'hDDD2313E2D1BAC08AC86DAC33D2E2391FCB133DCD7262BEA38796DBD728F11EF),
.INIT_10(256'h031A330008006900C61E5A00C9000000E1040000AE0000004D00000006000000),
.INIT_11(256'h3E34F700272EBF00E6FB4800FBE5000039CFC40064CBD60088001200D1000000),
.INIT_12(256'h8B9669000C0033004E920000CD005A0033880000F00000009F8C000058000000),
.INIT_13(256'h1E9790BA18924B2979E790057BE64B96D5FA6F2C97E1EEBFDB8A06939D958700),
.INIT_14(256'h55AB69DD770E1A62B799CC002E870000525038BF34EB1100BB00960066000000),
.INIT_15(256'h1BF6DEAE2B53BF11977CDE001C620000F9E88FCC8D53B4737E008400B1000000),
.INIT_16(256'h89BFFFDD27968C626B8D5A007E1F9600D444F4BF3E73DD003D145A006C98CC00),
.INIT_17(256'h0DAF17762215E55A3E9AA867AA9BE5F423278A82488322AE1B703EF1CB6F2962),
.INIT_18(256'hF8E1C8FBF3FB92FB3DE5A1FB32FBFBFB1AFFFBFB55FBFBFBB6FBFBFBFDFBFBFB),
.INIT_19(256'hC5CF0CFBDCD544FB1D00B3FB001EFBFBC2343FFB9F302DFB73FBE9FB2AFBFBFB),
.INIT_1A(256'h706D92FBF7FBC8FBB569FBFB36FBA1FBC873FBFB0BFBFBFB6477FBFBA3FBFBFB),
.INIT_1B(256'hE56C6B41E369B0D2821C6BFE801DB06D2E0194D76C1A15442071FD68666E7CFB),
.INIT_1C(256'hAE5092268CF5E1994C6237FBD57CFBFBA9ABC344CF10EAFB40FB6DFB9DFBFBFB),
.INIT_1D(256'hE00D2555D0A844EA6C8725FBE799FBFB0213743776A84F8885FB7FFB4AFBFBFB),
.INIT_1E(256'h72440426DC6D77999076A1FB85E46DFB2FBF0F44C58826FBC6EFA1FB976337FB),
.INIT_1F(256'hF654EC8DD9EE1EA1C561539C51601E0FD8DC7179B378D955E08BC50A3094D299),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
