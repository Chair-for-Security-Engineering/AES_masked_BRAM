//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_1_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hF8185D8EC6C3665000000000000000002BE2F40E2A06F0EF0000000000000000),
.INIT_01(256'hE54E72D8F852248FA91F77F3ECBE7C1C80AF745A735DCCE3150ED2FB817E08C5),
.INIT_02(256'hCC3DE4C47610FF4824B62959FF1F565470E4F0B5E4E7C517F72928143D914608),
.INIT_03(256'h85D9902F4E61B4782DEFF1E3E1B5D753F1655522C5228E8A3C1F2BD83085CDA8),
.INIT_04(256'hF5410DA49D06CA4C1A8C07BF28749FED2D4E6917A9E542138DE556106CCE1D91),
.INIT_05(256'h73C00995D9A14215EB8798E87D3FEAB4D1180EE8464478550C33A0839889D0DD),
.INIT_06(256'hD568CF8D78986976180467B7B014C1A9DBFDAF768BF0F470E54B8EEC8F99EA30),
.INIT_07(256'h134F84152ECBFCD45D5D43BD035F5DFF1973F95E08DBADB3AEB1BD5CE3A0B00D),
.INIT_08(256'h05E5A0733B3E9BADFDFDFDFDFDFDFDFDD61F09F3D7FB0D12FDFDFDFDFDFDFDFD),
.INIT_09(256'h18B38F2505AFD97254E28A0E114381E17D5289A78EA0311EE8F32F067C83F538),
.INIT_0A(256'h31C019398BED02B5D94BD4A402E2ABA98D190D48191A38EA0AD4D5E9C06CBBF5),
.INIT_0B(256'h78246DD2B39C4985D0120C1E1C482AAE0C98A8DF38DF7377C1E2D625CD783055),
.INIT_0C(256'h08BCF05960FB37B1E771FA42D5896210D0B394EA5418BFEE7018ABED9133E06C),
.INIT_0D(256'h8E3DF468245CBFE8167A651580C217492CE5F315BBB985A8F1CE5D7E65742D20),
.INIT_0E(256'h289532708565948BE5F99A4A4DE93C542600528B760D098D18B67311726417CD),
.INIT_0F(256'hEEB279E8D3360129A0A0BE40FEA2A002E48E04A3F526504E534C40A11E5D4DF0),
.INIT_10(256'h57EEBEAFDABF37FA0000000000000000C2121C64505C8A2E0000000000000000),
.INIT_11(256'h5EDF01FF16595F6FB658CBF27C801338ECB76145E2777993CE9356DC5D12D74F),
.INIT_12(256'h01C9F2CCDF11A49C47CCD401FFAEE0EFE01B9C91926F666D76A75DD27D76DA8F),
.INIT_13(256'h6116B1E7E98AA3E127C55C37C6EC238031C68B5D4CAF6CAEF8F3DE5CF3304B01),
.INIT_14(256'hF4491267B2450C330D18E99C79FAC1229062C6FCBD05B3C39EADFDAE9E3BA164),
.INIT_15(256'h7A9C10E93C821CBD4FD7ECC33428D9726C765356185A6D30F1FC308AA72E2816),
.INIT_16(256'h2B2B4FD97BEBCBCDC3912C404A5475559580F97A1D98A5B6CFE11F0F81E381DD),
.INIT_17(256'hAE72D34E6D33D6C9356D08B92026DF30F48E645FB64EE0598215651B09C02C0C),
.INIT_18(256'hAA1343522742CA07FDFDFDFDFDFDFDFD3FEFE199ADA177D3FDFDFDFDFDFDFDFD),
.INIT_19(256'hA322FC02EBA4A2924BA5360F817DEEC5114A9CB81F8A846E336EAB21A0EF2AB2),
.INIT_1A(256'hFC340F3122EC5961BA3129FC02531D121DE6616C6F929B908B5AA02F808B2772),
.INIT_1B(256'h9CEB4C1A14775E1CDA38A1CA3B11DE7DCC3B76A0B1529153050E23A10ECDB6FC),
.INIT_1C(256'h09B4EF9A4FB8F1CEF0E5146184073CDF6D9F3B0140F84E3E6350005363C65C99),
.INIT_1D(256'h8761ED14C17FE140B22A113EC9D5248F918BAEABE5A790CD0C01CD775AD3D5EB),
.INIT_1E(256'hD6D6B224861636303E6CD1BDB7A988A8687D0487E065584B321CE2F27C1E7C20),
.INIT_1F(256'h538F2EB390CE2B34C890F544DDDB22CD097399A24BB31DA47FE898E6F43DD1F1),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
