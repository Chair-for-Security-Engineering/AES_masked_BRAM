//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_7_x26_x49(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'h2D61703FA9003800F25E9C00AC000E004C00ED002C001F008500170000000000),
.INIT_01(256'hBDBAD2E40C0AAF0A958FC9D1FE006E00AA0039002E002F009E003E00FF00CD00),
.INIT_02(256'h4E1371CDF63C05BC714FFD114C000C00CEDF0D5F8380D2005B002B00AC004E00),
.INIT_03(256'h6A9A6744B53674B6A2CC1C92F8008A009C8D6D0D67800400F452B652B5006500),
.INIT_04(256'hCED6BD8837008800B78DF7D3F0007C0082640D644C005100ED005100A2008C00),
.INIT_05(256'h8F907E7EA2769FC601C1C32F927C9CCC79357485B2B02D00EB51D5E1A1B00D00),
.INIT_06(256'h0C1D1DC3C98514059525377BB1B9DFB918BBF53BFB8084002B0075001600DA00),
.INIT_07(256'hF9096A67BAF3E5C3973BB7D535C5D97557B83888E3301E00990345B3F3B0BD00),
.INIT_08(256'hD09C8DC254FDC5FD0FA361FD51FDF3FDB1FD10FDD1FDE2FD78FDEAFDFDFDFDFD),
.INIT_09(256'h40472F19F1F752F76872342C03FD93FD57FDC4FDD3FDD2FD63FDC3FD02FD30FD),
.INIT_0A(256'hB3EE8C300BC1F8418CB200ECB1FDF1FD3322F0A27E7D2FFDA6FDD6FD51FDB3FD),
.INIT_0B(256'h97679AB948CB894B5F31E16F05FD77FD617090F09A7DF9FD09AF4BAF48FD98FD),
.INIT_0C(256'h332B4075CAFD75FD4A700A2E0DFD81FD7F99F099B1FDACFD10FDACFD5FFD71FD),
.INIT_0D(256'h726D83835F8B623BFC3C3ED26F81613184C889784F4DD0FD16AC281C5C4DF0FD),
.INIT_0E(256'hF1E0E03E3478E9F868D8CA864C442244E54608C6067D79FDD6FD88FDEBFD27FD),
.INIT_0F(256'h04F4979A470E183E6AC64A28C8382488AA45C5751ECDE3FD64FEB84E0E4D40FD),
.INIT_10(256'hB332579265003F0041A010003300DC00AB0000005E00EB00C300DD0000000000),
.INIT_11(256'h34A3C20383F2CBF21FC35C630C00F1005800E100AF0008001B001700DA00C800),
.INIT_12(256'h0994B4B4824781C794CC1C6C36000000270DD58DE3800F00E700200098004100),
.INIT_13(256'h4435EB159EB58F35009F9A3FF300D7001E3DFEBDE8801600F5302030B8007300),
.INIT_14(256'h8F658FC580003E00E2D6577668006300B021FF21EA00BB004700BD000A00EE00),
.INIT_15(256'h6CDE1919BE647503D89F18588F96F1F1D6FAEC9D326716000ADB85BCF9676800),
.INIT_16(256'hDEFB87DB8C7F6BFFDC82B02286385438EF2CF9AC84808C00B000930041007C00),
.INIT_17(256'hF770DB37481BDAFC2CFB353C9BAE3CC943C72020A6E7DB0037EB618C48670000),
.INIT_18(256'h4ECFAA6F98FDC2FDBC5DEDFDCEFD21FD56FDFDFDA3FD16FD3EFD20FDFDFDFDFD),
.INIT_19(256'hC95E3FFE7E0F360FE23EA19EF1FD0CFDA5FD1CFD52FDF5FDE6FDEAFD27FD35FD),
.INIT_1A(256'hF46949497FBA7C3A6931E191CBFDFDFDDAF028701E7DF2FD1AFDDDFD65FDBCFD),
.INIT_1B(256'hB9C816E8634872C8FD6267C20EFD2AFDE3C00340157DEBFD08CDDDCD45FD8EFD),
.INIT_1C(256'h729872387DFDC3FD1F2BAA8B95FD9EFD4DDC02DC17FD46FDBAFD40FDF7FD13FD),
.INIT_1D(256'h9123E4E4439988FE2562E5A5726B0C0C2B071160CF9AEBFDF7267841049A95FD),
.INIT_1E(256'h23067A2671829602217F4DDF7BC5A9C512D10451797D71FD4DFD6EFDBCFD81FD),
.INIT_1F(256'h0A8D26CAB5E62701D106C8C16653C134BE3ADDDD5B1A26FDCA169C71B59AFDFD),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
