//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_7_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'h2D61703FA9003800F25E9C00AC000E004C00ED002C001F008500170000000000),
.INIT_01(256'hBDBAD2E40C0AAF0A958FC9D1FE006E00AA0039002E002F009E003E00FF00CD00),
.INIT_02(256'h4E1371CDF63C05BC714FFD114C000C00CEDF0D5F8380D2005B002B00AC004E00),
.INIT_03(256'h6A9A6744B53674B6A2CC1C92F8008A009C8D6D0D67800400F452B652B5006500),
.INIT_04(256'hCED6BD8837008800B78DF7D3F0007C0082640D644C005100ED005100A2008C00),
.INIT_05(256'h8F907E7EA2769FC601C1C32F927C9CCC79357485B2B02D00EB51D5E1A1B00D00),
.INIT_06(256'h0C1D1DC3C98514059525377BB1B9DFB918BBF53BFB8084002B0075001600DA00),
.INIT_07(256'hF9096A67BAF3E5C3973BB7D535C5D97557B83888E3301E00990345B3F3B0BD00),
.INIT_08(256'hD09C8DC254FDC5FD0FA361FD51FDF3FDB1FD10FDD1FDE2FD78FDEAFDFDFDFDFD),
.INIT_09(256'h40472F19F1F752F76872342C03FD93FD57FDC4FDD3FDD2FD63FDC3FD02FD30FD),
.INIT_0A(256'hB3EE8C300BC1F8418CB200ECB1FDF1FD3322F0A27E7D2FFDA6FDD6FD51FDB3FD),
.INIT_0B(256'h97679AB948CB894B5F31E16F05FD77FD617090F09A7DF9FD09AF4BAF48FD98FD),
.INIT_0C(256'h332B4075CAFD75FD4A700A2E0DFD81FD7F99F099B1FDACFD10FDACFD5FFD71FD),
.INIT_0D(256'h726D83835F8B623BFC3C3ED26F81613184C889784F4DD0FD16AC281C5C4DF0FD),
.INIT_0E(256'hF1E0E03E3478E9F868D8CA864C442244E54608C6067D79FDD6FD88FDEBFD27FD),
.INIT_0F(256'h04F4979A470E183E6AC64A28C8382488AA45C5751ECDE3FD64FEB84E0E4D40FD),
.INIT_10(256'h9501A71F8C00EB00331EA900E90026004E00AD000C00A4009E00D50000000000),
.INIT_11(256'hAB074E19F95F495F8447C95915000D00C500F1009500EA00C3005F004F009800),
.INIT_12(256'h70959502EBCC5B450BADCFB3B8002900076233EB74890B004F005A000B005500),
.INIT_13(256'h5A00689719937E1AA867BB79C300850098F17B786A89C2000693C493C3004A00),
.INIT_14(256'h5ACA08D41E001900526AA8746A00C500D3BF50BFB8007000AD008600A500C500),
.INIT_15(256'hAD66124267308D0A2C993BBD9A6FD855C440AA7A783A5D006CFFAAC5B33A3E00),
.INIT_16(256'hDDF058671B62CBEB0877AC6959AEA8AE56DD02540C891300B000C50062005C00),
.INIT_17(256'h3ECF5662E552D8E162172B332EC132FB55B1EC024BB3B900656CFD56F33A2000),
.INIT_18(256'h68FC5AE271FD16FDCEE354FD14FDDBFDB3FD50FDF1FD59FD63FD28FDFDFDFDFD),
.INIT_19(256'h56FAB3E404A2B4A279BA34A4E8FDF0FD38FD0CFD68FD17FD3EFDA2FDB2FD65FD),
.INIT_1A(256'h8D6868FF1631A6B8F650324E45FDD4FDFA9FCE168974F6FDB2FDA7FDF6FDA8FD),
.INIT_1B(256'hA7FD956AE46E83E7559A46843EFD78FD650C868597743FFDFB6E396E3EFDB7FD),
.INIT_1C(256'hA737F529E3FDE4FDAF97558997FD38FD2E42AD4245FD8DFD50FD7BFD58FD38FD),
.INIT_1D(256'h509BEFBF9ACD70F7D164C640679225A839BD578785C7A0FD910257384EC7C3FD),
.INIT_1E(256'h200DA59AE69F3616F58A5194A4535553AB20FFA9F174EEFD4DFD38FD9FFDA1FD),
.INIT_1F(256'hC332AB9F18AF251C9FEAD6CED33CCF06A84C11FFB64E44FD989100AB0EC7DDFD),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
