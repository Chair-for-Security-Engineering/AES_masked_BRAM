//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_1_x26_x49(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hF8185D8EC6C3665000000000000000002BE2F40E2A06F0EF0000000000000000),
.INIT_01(256'hE54E72D8F852248FA91F77F3ECBE7C1C80AF745A735DCCE3150ED2FB817E08C5),
.INIT_02(256'hCC3DE4C47610FF4824B62959FF1F565470E4F0B5E4E7C517F72928143D914608),
.INIT_03(256'h85D9902F4E61B4782DEFF1E3E1B5D753F1655522C5228E8A3C1F2BD83085CDA8),
.INIT_04(256'hF5410DA49D06CA4C1A8C07BF28749FED2D4E6917A9E542138DE556106CCE1D91),
.INIT_05(256'h73C00995D9A14215EB8798E87D3FEAB4D1180EE8464478550C33A0839889D0DD),
.INIT_06(256'hD568CF8D78986976180467B7B014C1A9DBFDAF768BF0F470E54B8EEC8F99EA30),
.INIT_07(256'h134F84152ECBFCD45D5D43BD035F5DFF1973F95E08DBADB3AEB1BD5CE3A0B00D),
.INIT_08(256'h05E5A0733B3E9BADFDFDFDFDFDFDFDFDD61F09F3D7FB0D12FDFDFDFDFDFDFDFD),
.INIT_09(256'h18B38F2505AFD97254E28A0E114381E17D5289A78EA0311EE8F32F067C83F538),
.INIT_0A(256'h31C019398BED02B5D94BD4A402E2ABA98D190D48191A38EA0AD4D5E9C06CBBF5),
.INIT_0B(256'h78246DD2B39C4985D0120C1E1C482AAE0C98A8DF38DF7377C1E2D625CD783055),
.INIT_0C(256'h08BCF05960FB37B1E771FA42D5896210D0B394EA5418BFEE7018ABED9133E06C),
.INIT_0D(256'h8E3DF468245CBFE8167A651580C217492CE5F315BBB985A8F1CE5D7E65742D20),
.INIT_0E(256'h289532708565948BE5F99A4A4DE93C542600528B760D098D18B67311726417CD),
.INIT_0F(256'hEEB279E8D3360129A0A0BE40FEA2A002E48E04A3F526504E534C40A11E5D4DF0),
.INIT_10(256'h2C4CB2679CCA48AB0000000000000000FA92E934D886816A0000000000000000),
.INIT_11(256'h1F69D405DE9C698CDDE0577884BB38150299DDE1329D9199E43CF73DDE04FB33),
.INIT_12(256'h0E72B5A531C744DE03BAA6C6010420FC8F6625A04E2D2A2593B7AA57FD654001),
.INIT_13(256'hF86839D7869EBFD995EB9520FE3E4C479575DC42761EC7D11B1D1ED37FC7C8BB),
.INIT_14(256'h1A11CD974AF96C8E70A5DBEAB1EAA11EE9BB17145DB752E936B23959818B35DB),
.INIT_15(256'hE4B7011179905BF17BDD3D6D5F7594482DC278D43762A5B3F5E78E6AC45A325A),
.INIT_16(256'hC80C84C8DC1CE5ADD96669EBD15C5EEE5454AD25C8CC44C83744BFF1256492EE),
.INIT_17(256'hA1C7F00C48285AA0CBFDB9A016106D4420675D8022631CC7CAD519296E41B4B4),
.INIT_18(256'hD1B14F9A6137B556FDFDFDFDFDFDFDFD076F14C9257B7C97FDFDFDFDFDFDFDFD),
.INIT_19(256'hE29429F823619471201DAA857946C5E8FF64201CCF606C6419C10AC023F906CE),
.INIT_1A(256'hF38F4858CC3AB923FE475B3BFCF9DD01729BD85DB3D0D7D86E4A57AA0098BDFC),
.INIT_1B(256'h0595C42A7B634224681668DD03C3B1BA688821BF8BE33A2CE6E0E32E823A3546),
.INIT_1C(256'hE7EC306AB70491738D5826174C175CE31446EAE9A04AAF14CB4FC4A47C76C826),
.INIT_1D(256'h194AFCEC846DA60C8620C090A28869B5D03F8529CA9F584E081A739739A7CFA7),
.INIT_1E(256'h35F1793521E11850249B94162CA1A313A9A950D83531B935CAB9420CD8996F13),
.INIT_1F(256'h5C3A0DF1B5D5A75D3600445DEBED90B9DD9AA07DDF9EE13A3728E4D493BC4949),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
