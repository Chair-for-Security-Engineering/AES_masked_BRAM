//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_2_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hA2C219493CB99CBB70DCB428D07C0A04543411E30000000055D0150200000000),
.INIT_01(256'h3EEA3EDA8356D6A158BDCB1EBDBC7EDD7E079972D82534C9C1A0CF3C00000000),
.INIT_02(256'h580695FB428B305B69FBDB7912F21A58C1D320A0000000009F687B1E00000000),
.INIT_03(256'h909CE9D5FB8473AEE1DC0B068D26939AC12C8DF2A0BB4358D52070178C6A8365),
.INIT_04(256'hC35554F20BB22D36069EAE0694C688783E56916BEF2DAF6DB4FB5E8300000000),
.INIT_05(256'hB1939D8FBB52682303D2FC1D35CA306D36473BD8F4CB5867C16A655C00000000),
.INIT_06(256'h2D9DA32320CDBBF43987880631379034060462F203D92CF6E1C4C077DEC6B1A9),
.INIT_07(256'h1FFD25F782D9E31A88996140763BC12E30CDF99674B5B8795E793E8B46B826D8),
.INIT_08(256'h5939E2B2C74267408B274FD32B87F1FFAFCFEA18FBFBFBFBAE2BEEF9FBFBFBFB),
.INIT_09(256'hC511C52178AD2D5AA34630E54647852685FC628923DECF323A5B34C7FBFBFBFB),
.INIT_0A(256'hA3FD6E00B970CBA092002082E909E1A33A28DB5BFBFBFBFB649380E5FBFBFBFB),
.INIT_0B(256'h6B67122E007F88551A27F0FD76DD68613AD776095B40B8A32EDB8BEC7791789E),
.INIT_0C(256'h38AEAF09F049D6CDFD6555FD6F3D7383C5AD6A9014D654964F00A578FBFBFBFB),
.INIT_0D(256'h4A68667440A993D8F82907E6CE31CB96CDBCC0230F30A39C3A919EA7FBFBFBFB),
.INIT_0E(256'hD66658D8DB36400FC27C73FDCACC6BCFFDFF9909F822D70D1A3F3B8C253D4A52),
.INIT_0F(256'hE406DE0C792218E173629ABB8DC03AD5CB36026D8F4E4382A582C570BD43DD23),
.INIT_10(256'hD74F2C30D656B4FBD0FD18B15CB5092F5311D4DD00000000C15F429700000000),
.INIT_11(256'h836C442F47A20B213BB7040C7D27CD5820A67EB3EF3924F252DEC30400000000),
.INIT_12(256'h435B8C1011CBCBDEEA47163FDE6D334FB32BB86B00000000CA8EC5CA00000000),
.INIT_13(256'h7E9618747A421BECD75C4946BA3D276F3FE478E883D2DD8C19C8910BD35446C1),
.INIT_14(256'hEAD3219C20972E5643DE5049BB7469699F5AAF2173629889C1C91E5D00000000),
.INIT_15(256'h5D13AA609745B7AA3804DC64CFB3F84B5A5BB3F9EF28CF08978D5A0B00000000),
.INIT_16(256'hF78290612B0A05EBF0214F1AF5AC0791588B7CE411CC62BFEDF3267362AEFA36),
.INIT_17(256'h4BCE858404C7919D3FC8E291A6CB2486009068B3830FAE229912D515D398DE95),
.INIT_18(256'h2CB4D7CB2DAD4F002B06E34AA74EF2D4A8EA2F26FBFBFBFB3AA4B96CFBFBFBFB),
.INIT_19(256'h7897BFD4BC59F0DAC04CFFF786DC36A3DB5D854814C2DF09A92538FFFBFBFBFB),
.INIT_1A(256'hB8A077EBEA30302511BCEDC42596C8B448D04390FBFBFBFB31753E31FBFBFBFB),
.INIT_1B(256'h856DE38F81B9E0172CA7B2BD41C6DC94C41F831378292677E2336AF028AFBD3A),
.INIT_1C(256'h1128DA67DB6CD5ADB825ABB2408F929264A154DA889963723A32E5A6FBFBFBFB),
.INIT_1D(256'hA6E8519B6CBE4C51C3FF279F344803B0A1A0480214D334F36C76A1F0FBFBFBFB),
.INIT_1E(256'h0C796B9AD0F1FE100BDAB4E10E57FC6AA370871FEA3799441608DD88995501CD),
.INIT_1F(256'hB0357E7FFF3C6A66C433196A5D30DF7DFB6B934878F455D962E92EEE2863256E),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
