//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_3_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
		.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hD21EAD61ECC596BF000000000000000001E404E1000000000000000000000000),
.INIT_01(256'h4E368AF2532ADCA528617F366DC074D92BD78C70D82534C99470DA3E00000000),
.INIT_02(256'h28DA21D392F73A5F19276F51C28E105C940335A200000000CAB86E1C00000000),
.INIT_03(256'hE0405DFD2BF879AA9100BF2E5D5A999E94FC98F0A0BB435880F065158C6A8365),
.INIT_04(256'hB389E0DADBCE273276421A2E44BA827C6B868469EF2DAF6DE12B4B8100000000),
.INIT_05(256'hC14F29A76B2E6227730E4835E5B63A6963972EDAF4CB586794BA705E00000000),
.INIT_06(256'h5D41170BF0B1B1F0495B3C2EE14B9A3053D477F003D92CF6B414D575DEC6B1A9),
.INIT_07(256'h6F2191DF52A5E91EF845D568A647CB2A651DEC9474B5B8790BA92B8946B826D8),
.INIT_08(256'h25E95A961B326148F7F7F7F7F7F7F7F7F613F316F7F7F7F7F7F7F7F7F7F7F7F7),
.INIT_09(256'hB9C17D05A4DD2B52DF9688C19A37832EDC207B872FD2C33E63872DC9F7F7F7F7),
.INIT_0A(256'hDF2DD6246500CDA8EED098A63579E7AB63F4C255F7F7F7F73D4F99EBF7F7F7F7),
.INIT_0B(256'h17B7AA0ADC0F8E5D66F748D9AAAD6E69630B6F07574CB4AF770792E27B9D7492),
.INIT_0C(256'h447E172D2C39D0C581B5EDD9B34D758B9C71739E18DA589A16DCBC76F7F7F7F7),
.INIT_0D(256'h36B8DE509CD995D084F9BFC21241CD9E9460D92D033CAF90634D87A9F7F7F7F7),
.INIT_0E(256'hAAB6E0FC07464607BEACCBD916BC6DC7A4238007F42EDB0143E322822931465E),
.INIT_0F(256'h98D66628A5521EE90FB2229F51B03CDD92EA1B6383424F8EFC5EDC7EB14FD12F),
.INIT_10(256'h07B234818AE3BDD40000000000000000924E964A000000000000000000000000),
.INIT_11(256'h53915C9E1B17020EEB4A1CBD2192C477E1F93C24EF3924F29381819300000000),
.INIT_12(256'h93A694A14D7EC2F13ABA0E8E82D83A607274FAFC000000000BD1875D00000000),
.INIT_13(256'hAE6B00C526F712C307A151F7E6882E40FEBB3A7F83D2DD8CD897D39CD35446C1),
.INIT_14(256'h3A2E392D7C222779932348F8E7C160465E05EDB67362988900965CCA00000000),
.INIT_15(256'h8DEEB2D1CBF0BE85E8F9C4D59306F1649B04F16EEF28CF0856D2189C00000000),
.INIT_16(256'h277F88D077BF0CC420DC57ABA9190EBE99D43E7311CC62BF2CAC64E462AEFA36),
.INIT_17(256'h9B339D35587298B2EF35FA20FA7E2DA9C1CF2A24830FAE22584D9782D398DE95),
.INIT_18(256'hF045C3767D144A23F7F7F7F7F7F7F7F765B961BDF7F7F7F7F7F7F7F7F7F7F7F7),
.INIT_19(256'hA466AB69ECE0F5F91CBDEB4AD6653380160ECBD318CED30564767664F7F7F7F7),
.INIT_1A(256'h64516356BA893506CD4DF979752FCD9785830D0BF7F7F7F7FC2670AAF7F7F7F7),
.INIT_1B(256'h599CF732D100E534F056A600117FD9B7094CCD8874252A7B2F60246B24A3B136),
.INIT_1C(256'hCDD9CEDA8BD5D08E64D4BF0F103697B1A9F21A4184956F7EF761AB3DF7F7F7F7),
.INIT_1D(256'h7A1945263C0749721F0E332264F106936CF3069918DF38FFA125EF6BF7F7F7F7),
.INIT_1E(256'hD0887F278048FB33D72BA05C5EEEF9496E23C984E63B9548DB5B931395590DC1),
.INIT_1F(256'h6CC46AC2AF856F4518C20DD70D89DA5E3638DDD374F859D5AFBA6075246F2962),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
