//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_9_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
		.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hAC7AE500497A00000000000000000000D600E500330000000000000000000000),
.INIT_01(256'h6CD8B500C7965000D14EAD009F00AD00BBA2180010ECFD007C4E000032000000),
.INIT_02(256'hEEA8970079A8000042D2720030D2000046009700D100000090007200E2000000),
.INIT_03(256'h1FDDF9D894C13C8A56BF152C38A3357E640B2AA6EF17EFF45713C652390FE600),
.INIT_04(256'hAC6821F887A6A09C7AAAFE00D000FE00B48E43649F40C20084AA00002E000000),
.INIT_05(256'hAF09B23BCA89335FABE453004F0053001AEF7DA77F6FFCC3F8E400001C000000),
.INIT_06(256'hABE779CAF2298AAE4F17940097BDE60061D31B56381DE83263C56A00BB6F1800),
.INIT_07(256'h8D45C0C5C89761F34F6EE7388BD8C76A940F7127D1DDD011B0C2CA467474EA14),
.INIT_08(256'h5B8D12F7BE8DF7F7F7F7F7F7F7F7F7F721F712F7C4F7F7F7F7F7F7F7F7F7F7F7),
.INIT_09(256'h9B2F42F73061A7F726B95AF768F75AF74C55EFF7E71B0AF78BB9F7F7C5F7F7F7),
.INIT_0A(256'h195F60F78E5FF7F7B52585F7C725F7F7B1F760F726F7F7F767F785F715F7F7F7),
.INIT_0B(256'hE82A0E2F6336CB7DA148E2DBCF54C28993FCDD5118E01803A0E431A5CEF811F7),
.INIT_0C(256'h5B9FD60F7051576B8D5D09F727F709F74379B49368B735F7735DF7F7D9F7F7F7),
.INIT_0D(256'h58FE45CC3D7EC4A85C13A4F7B8F7A4F7ED188A5088980B340F13F7F7EBF7F7F7),
.INIT_0E(256'h5C108E3D05DE7D59B8E063F7604A11F79624ECA1CFEA1FC594329DF74C98EFF7),
.INIT_0F(256'h7AB237323F609604B89910CF7C2F309D63F886D0262A27E647353DB183831DE3),
.INIT_10(256'h4337DC009F37000000000000000000007400DC00A80000000000000000000000),
.INIT_11(256'h28EEB900E6FC65007612B3006400B300ACD90A0062CBD600C5120000D7000000),
.INIT_12(256'h7F8F0600798F00003CB8DA00E6B80000F0000600F60000008400DA005E000000),
.INIT_13(256'hBC795EBA3BF8CB295D3AEB0506BBA29616607B2C91E1EEBFC014CE939B958700),
.INIT_14(256'h7E5D36DD41BE55621A5C2600460026000D0872BF32EB11003C5C000060000000),
.INIT_15(256'h66F720AE4B0643116C4E950022009500A6A2D7CC8B53B473F94E0000B7000000),
.INIT_16(256'h167D20DDF39E9962727C3000F420EA00DD9064BF3873DD00ECC416006A98CC00),
.INIT_17(256'hC49A6976A0F8435A719C636776412AF42AE108824E8322AECAB260F1CD6F2962),
.INIT_18(256'hB4C02BF768C0F7F7F7F7F7F7F7F7F7F783F72BF75FF7F7F7F7F7F7F7F7F7F7F7),
.INIT_19(256'hDF194EF7110B92F781E544F793F744F75B2EFDF7953C21F732E5F7F720F7F7F7),
.INIT_1A(256'h8878F1F78E78F7F7CB4F2DF7114FF7F707F7F1F701F7F7F773F72DF7A9F7F7F7),
.INIT_1B(256'h4B8EA94DCC0F3CDEAACD1CF2F14C5561E1978CDB6616194837E339646C6270F7),
.INIT_1C(256'h89AAC12AB649A295EDABD1F7B1F7D1F7FAFF8548C51CE6F7CBABF7F797F7F7F7),
.INIT_1D(256'h9100D759BCF1B4E69BB962F7D5F762F75155203B7CA443840EB9F7F740F7F7F7),
.INIT_1E(256'hE18AD72A04696E95858BC7F703D71DF72A679348CF842AF71B33E1F79D6F3BF7),
.INIT_1F(256'h336D9E81570FB4AD866B949081B6DD03DD16FF75B974D5593D4597063A98DE95),


	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
