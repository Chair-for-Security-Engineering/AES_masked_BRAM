//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_4_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
		.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hF28994117D1100006820AB2EDD82000098C40000DD1300004728000007FA0000),
.INIT_01(256'h773E23A6015F0000671D7AFF4D200000D5BB6666B844000080DD00008E410000),
.INIT_02(256'hFEE415139B96CF4C74DEBA3F74C90000EBD62CAF55FA73F0981500007C630000),
.INIT_03(256'hFED6282E625D45C60A921590951A7E7E5D52BE3DCB56870450EF0000FAD70000),
.INIT_04(256'hE0B5DB5E16549C9CA6C078FD6A1B000003710000EC0C00009CDD000076A50000),
.INIT_05(256'hFED5478E102C561AF1E94188434C0945191581CD3FA1064ACFF024688A27C589),
.INIT_06(256'hF0C4292FAD8E61E2941028ADAC3F00006C7F5FDC39B841C26DCE414162530000),
.INIT_07(256'h7F352B613A6735FAA65C7BB2E00D632F99F43EF105FAA76825F8713D85CAD19D),
.INIT_08(256'h1D667BFE92FEEFEF87CF44C1326DEFEF772BEFEF32FCEFEFA8C7EFEFE815EFEF),
.INIT_09(256'h98D1CC49EEB0EFEF88F29510A2CFEFEF3A54898957ABEFEF6F32EFEF61AEEFEF),
.INIT_0A(256'h110BFAFC747920A39B3155D09B26EFEF0439C340BA159C1F77FAEFEF938CEFEF),
.INIT_0B(256'h1139C7C18DB2AA29E57DFA7F7AF59191B2BD51D224B968EBBF00EFEF1538EFEF),
.INIT_0C(256'h0F5A34B1F9BB7373492F971285F4EFEFEC9EEFEF03E3EFEF7332EFEF994AEFEF),
.INIT_0D(256'h113AA861FFC3B9F51E06AE67ACA3E6AAF6FA6E22D04EE9A5201FCB8765C82A66),
.INIT_0E(256'h1F2BC6C042618E0D7BFFC74243D0EFEF8390B033D657AE2D8221AEAE8DBCEFEF),
.INIT_0F(256'h90DAC48ED588DA1549B3945D0FE28CC0761BD11EEA154887CA179ED26A253E72),
.INIT_10(256'hBFCF4C166A0B000049915309874E00008F6A000008A60000511C0000D2D40000),
.INIT_11(256'h5FF81A40CE7800006D620A50E8F60000D3E10F0F49300000C953000058890000),
.INIT_12(256'h8E5A67C78F4A738969EFE0BA980F0000F0B1DD27101A36CC7A690000752D0000),
.INIT_13(256'hD2D118B897855AA04E1F2F75F4B4969686106D977BA6897377B300006AE50000),
.INIT_14(256'hA6B65A005B5A6262D961277D3F96000007820000DC120000321F0000ED8B0000),
.INIT_15(256'hC165B188BD081A790905B089617C0B6889B8E7848AF02D4E0B929BF803D15E3D),
.INIT_16(256'h4AFE3494268311EB24C2D18BB84F0000A58498625C3636CCC4B74545D2EA0000),
.INIT_17(256'hF3F394571E0F22BB95C7B28B87C4FF9C63F6A23B429CC65F0ACDBCDFCB473C5F),
.INIT_18(256'h5020A3F985E4EFEFA67EBCE668A1EFEF6085EFEFE749EFEFBEF3EFEF3D3BEFEF),
.INIT_19(256'hB017F5AF2197EFEF828DE5BF0719EFEF3C0EE0E0A6DFEFEF26BCEFEFB766EFEF),
.INIT_1A(256'h61B5882860A59C6686000F5577E0EFEF1F5E32C8FFF5D9239586EFEF9AC2EFEF),
.INIT_1B(256'h3D3EF757786AB54FA1F0C09A1B5B797969FF82789449669C985CEFEF850AEFEF),
.INIT_1C(256'h4959B5EFB4B58D8D368EC892D079EFEFE86DEFEF33FDEFEFDDF0EFEF0264EFEF),
.INIT_1D(256'h2E8A5E6752E7F596E6EA5F668E93E4876657086B651FC2A1E47D7417EC3EB1D2),
.INIT_1E(256'hA511DB7BC96CFE04CB2D3E6457A0EFEF4A6B778DB3D9D9232B58AAAA3D05EFEF),
.INIT_1F(256'h1C1C7BB8F1E0CD547A285D64682B10738C194DD4AD7329B0E522533024A8D3B0),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
