//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_0_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'h8E3EE8A610456D547626B528D6860B0478C8E00C2CFCF1EF532A140206FA0100),
.INIT_01(256'h9368C7F02ED42F8BDF39C2DB3A387718D385605875A7CDE34624C6F9878409C5),
.INIT_02(256'hBA1B51ECA096F44C52909C7129995D5023CEE4B7E21DC417A4033C163B6B4708),
.INIT_03(256'hF3FF250798E7BF7C5BC944CB3733DC57A24F4120C3D88F8A6F353FDA367FCCA8),
.INIT_04(256'h8367B88C4B80C1486CAAB297FEF294E97E647D15AF1F4313DECF42126A341C91),
.INIT_05(256'h05E6BCBD0F2749119DA12DC0ABB9E1B082321AEA40BE79555F19B4819E73D1DD),
.INIT_06(256'hA34E7AA5AE1E62726E22D29F6692CAAD88D7BB748D0AF570B6619AEE8963EB30),
.INIT_07(256'h6569313DF84DF7D02B7BF695D5D956FB4A59ED5C0E21ACB3FD9BA95EE55AB10D),
.INIT_08(256'h70C01658EEBB93AA88D84BD62878F5FA86361EF2D2020F11ADD4EAFCF804FFFE),
.INIT_09(256'h6D96390ED02AD17521C73C25C4C689E62D7B9EA68B59331DB8DA3807797AF73B),
.INIT_0A(256'h44E5AF125E680AB2AC6E628FD767A3AEDD301A491CE33AE95AFDC2E8C595B9F6),
.INIT_0B(256'h0D01DBF966194182A537BA35C9CD22A95CB1BFDE3D26717491CBC124C8813256),
.INIT_0C(256'h7D994672B57E3FB692544C69000C6A17809A83EB51E1BDED2031BCEC94CAE26F),
.INIT_0D(256'hFB184243F1D9B7EF635FD33E55471F4E7CCCE414BE4087ABA1E74A7F608D2F23),
.INIT_0E(256'h5DB0845B50E09C8C90DC2C61986C34537629458A73F40B8E489F6410779D15CE),
.INIT_0F(256'h9B97CFC306B3092ED585086B2B27A805B4A713A2F0DF524D036557A01BA44FF3),
.INIT_10(256'h7490874975891F82237E39E6AF362878F0CE7FA4A3DFAB7932DC63C0F3832157),
.INIT_11(256'h7DA13819B96F77179526F214D3B63B40DE6B028511F458C4FC4F351CAE91F618),
.INIT_12(256'h22B7CB2A70278CE464B2EDE75098C897D2C7FF5161EC473A447B3E128EF5FBD8),
.INIT_13(256'h4268880146BC8B9904BB65D169DA0BF8031AE89DBF2C4DF9CA2FBD9C00B36A56),
.INIT_14(256'hD7372B811D73244B2E66D07AD6CCE95AA2BEA53C4E869294AC719E6E6DB88033),
.INIT_15(256'h59E2290F93B434C56CA9D5259B1EF10A5EAA3096EBD94C67C320534A54AD0941),
.INIT_16(256'h0855763FD4DDE3B5E0EF15A6E5625D2DA75C9ABAEE1B84E1FD3D7CCF7260A08A),
.INIT_17(256'h8D0CEAA8C205FEB11613315F8F10F748C652079F45CDC10EB0C906DBFA430D5B),
.INIT_18(256'h8A6E79B78B77E17CDD80C71851C8D6860E30815A5D215587CC229D3E0D7DDFA9),
.INIT_19(256'h835FC6E7479189E96BD80CEA2D48C5BE2095FC7BEF0AA63A02B1CBE2506F08E6),
.INIT_1A(256'hDC4935D48ED9721A9A4C1319AE6636692C3901AF9F12B9C4BA85C0EC700B0526),
.INIT_1B(256'hBC9676FFB8427567FA459B2F9724F506FDE4166341D2B30734D14362FE4D94A8),
.INIT_1C(256'h29C9D57FE38DDAB5D0982E84283217A45C405BC2B0786C6A528F609093467ECD),
.INIT_1D(256'hA71CD7F16D4ACA3B92572BDB65E00FF4A054CE681527B2993DDEADB4AA53F7BF),
.INIT_1E(256'hF6AB88C12A231D4B1E11EB581B9CA3D359A2644410E57A1F03C382318C9E5E74),
.INIT_1F(256'h73F214563CFB004FE8EDCFA171EE09B638ACF961BB333FF04E37F82504BDF3A5),

	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
	.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
