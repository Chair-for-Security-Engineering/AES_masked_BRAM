//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_6_x26(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hD161713F550039000E5E9D0050000F00B000EC00D0001E0079001600FC000100),
.INIT_01(256'h2DD6BF88FA00A400698FC8D102006F0030665E66D2002E0062003F000300CC00),
.INIT_02(256'hB21370CD0A3C04BC8D4FFC11B0000D0032DF0C5F7F80D300A7002A0050004F00),
.INIT_03(256'hD6DA26043D4201C272E031BE7A7EF57E54B958399B8005005A00E50049006400),
.INIT_04(256'hCA2E4470579C159C4B8DF6D30C007D001A006800B0005000110050005E008D00),
.INIT_05(256'hE704EBEAC8E00850FDC1C22F6E7C9DCC873777874EB02C001751D4E15DB00C00),
.INIT_06(256'hF01D1CC310A0302091DDCE83F4006700C19ED11E0780850096413541EA00DB00),
.INIT_07(256'h45492B2717A2B592BFEF62010E021FB2BAA928991F301F00761057A00FB0BC00),
.INIT_08(256'h2F9F8FC1ABFEC7FEF0A063FEAEFEF1FE4EFE12FE2EFEE0FE87FEE8FE02FEFFFE),
.INIT_09(256'hD328417604FE5AFE9771362FFCFE91FECE98A0982CFED0FE9CFEC1FEFDFE32FE),
.INIT_0A(256'h4CED8E33F4C2FA4273B102EF4EFEF3FECC21F2A1817E2DFE59FED4FEAEFEB1FE),
.INIT_0B(256'h2824D8FAC3BCFF3C8C1ECF4084800B80AA47A6C7657EFBFEA4FE1BFEB7FE9AFE),
.INIT_0C(256'h34D0BA8EA962EB62B573082DF2FE83FEE4FE96FE4EFEAEFEEFFEAEFEA0FE73FE),
.INIT_0D(256'h19FA1514361EF6AE033F3CD19082633279C98979B04ED2FEE9AF2A1FA34EF2FE),
.INIT_0E(256'h0EE3E23DEE5ECEDE6F23307D0AFE99FE3F602FE0F97E7BFE68BFCBBF14FE25FE),
.INIT_0F(256'hBBB7D5D9E95C4B6C41119CFFF0FCE14C4457D667E1CEE1FE88EEA95EF14E42FE),
.INIT_10(256'hE501D11FFC009D00431EDF00990050003E00DB007C00D200EE00A30070007600),
.INIT_11(256'h8B576849D6006000F447BF5965007B00BA0F880FE5009C00B30029003F00EE00),
.INIT_12(256'h0095E3029BCC2D457BADB9B3C8005F00776245EB04897D003F002C007B002300),
.INIT_13(256'h7F554BC2A05AC1D3DD62C87C25966596746D91E41A89B400E5002100B3003C00),
.INIT_14(256'hF717A3090C620D62226ADE741A00B3001C009900C8000600DD00F000D500B300),
.INIT_15(256'h50EBE9CF2A0DC6375C994DBDEA6FAE5504F06CCA083A2B001CFFDCC5C33A4800),
.INIT_16(256'h9BC61851A7AE7127939C318287007000DC278EAE7C8965008545F64512002A00),
.INIT_17(256'h2DAC43019057ABE4FCF9B3DD66F97CC343D7FC643BB3CF00C3BA5D80833A5600),
.INIT_18(256'h1BFF2FE102FE63FEBDE021FE67FEAEFEC0FE25FE82FE2CFE10FE5DFE8EFE88FE),
.INIT_19(256'h75A996B728FE9EFE0AB941A79BFE85FE44F176F11BFE62FE4DFED7FEC1FE10FE),
.INIT_1A(256'hFE6B1DFC6532D3BB8553474D36FEA1FE899CBB15FA7783FEC1FED2FE85FEDDFE),
.INIT_1B(256'h81ABB53C5EA43F2D239C3682DB689B688A936F1AE4774AFE1BFEDFFE4DFEC2FE),
.INIT_1C(256'h09E95DF7F29CF39CDC94208AE4FE4DFEE2FE67FE36FEF8FE23FE0EFE2BFE4DFE),
.INIT_1D(256'hAE151731D4F338C9A267B343149150ABFA0E9234F6C4D5FEE201223B3DC4B6FE),
.INIT_1E(256'h6538E6AF59508FD96D62CF7C79FE8EFE22D9705082779BFE7BBB08BBECFED4FE),
.INIT_1F(256'hD352BDFF6EA9551A02074D239807823DBD29029AC54D31FE3D44A37E7DC4A8FE),


	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
	.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
