//-----------------------------------------------------------------
//-- COMPANY : Ruhr University Bochum
//-- AUTHOR  : Aein Rezaei Shahmirzadi (aein.rezaeishahmirzadi@rub.de) and Amir Moradi (amir.moradi@rub.de) 
//-- DOCUMENT: [New First-Order Secure AES Performance Records](IACR Transactions on Cryptographic Hardware and Embeded Systems 2021(2))
//-- -----------------------------------------------------------------
//--
//-- Copyright (c) 2021, Aein Rezaei Shahmirzadi, Amir Moradi, 
//--
//-- All rights reserved.
//--
//-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
//-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
//-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
//-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
//-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
//-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
//-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
//-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//--
//-- Please see LICENSE and README for license and further instructions.
//--

module BRAM_2_x26_x49(
    input [9:0] ADDRA,
    input [9:0] ADDRB,
    input clk,
    input rst, input EN,
    output [7:0] DOA,
    output [7:0] DOB
    );



// Spartan-6
// Xilinx HDL Libraries Guide, version 14.7
//////////////////////////////////////////////////////////////////////////
// DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
// ===============|===========|===========|===============|=============//
// 19-36 | "18Kb" | 512 | 9-bit | 4-bit //
// 10-18 | "18Kb" | 1024 | 10-bit | 2-bit //
// 10-18 | "9Kb" | 512 | 9-bit | 2-bit //
// 5-9 | "18Kb" | 2048 | 11-bit | 1-bit //
// 5-9 | "9Kb" | 1024 | 10-bit | 1-bit //
// 3-4 | "18Kb" | 4096 | 12-bit | 1-bit //
// 3-4 | "9Kb" | 2048 | 11-bit | 1-bit //
// 2 | "18Kb" | 8192 | 13-bit | 1-bit //
// 2 | "9Kb" | 4096 | 12-bit | 1-bit //
// 1 | "18Kb" | 16384 | 14-bit | 1-bit //
// 1 | "9Kb" | 8192 | 12-bit | 1-bit //
//////////////////////////////////////////////////////////////////////////
BRAM_TDP_MACRO #(
	.BRAM_SIZE("9Kb"), // Target BRAM: "9Kb" or "18Kb"
	.DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6"
	.DOA_REG(1), // Optional port A output register (0 or 1)
	.DOB_REG(1), // Optional port B output register (0 or 1)
	.INIT_A(36'h0123), // Initial values on port A output port
	.INIT_B(36'h3210), // Initial values on port B output port
	.INIT_FILE ("NONE"),
	.READ_WIDTH_A (8), // Valid values are 1-36
	.READ_WIDTH_B (8), // Valid values are 1-36
	.SIM_COLLISION_CHECK ("NONE"), // Collision check enable "ALL", "WARNING_ONLY",
	// "GENERATE_X_ONLY" or "NONE"
	.SRVAL_A(36'h00000000), // Set/Reset value for port A output
	.SRVAL_B(36'h00000000), // Set/Reset value for port B output
	.WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
	.WRITE_WIDTH_A(8), // Valid values are 1-36
	.WRITE_WIDTH_B(8), // Valid values are 1-36
	
.INIT_00(256'hA2C219493CB99CBB70DCB428D07C0A04543411E30000000055D0150200000000),
.INIT_01(256'h3EEA3EDA8356D6A158BDCB1EBDBC7EDD7E079972D82534C9C1A0CF3C00000000),
.INIT_02(256'h580695FB428B305B69FBDB7912F21A58C1D320A0000000009F687B1E00000000),
.INIT_03(256'h909CE9D5FB8473AEE1DC0B068D26939AC12C8DF2A0BB4358D52070178C6A8365),
.INIT_04(256'hC35554F20BB22D36069EAE0694C688783E56916BEF2DAF6DB4FB5E8300000000),
.INIT_05(256'hB1939D8FBB52682303D2FC1D35CA306D36473BD8F4CB5867C16A655C00000000),
.INIT_06(256'h2D9DA32320CDBBF43987880631379034060462F203D92CF6E1C4C077DEC6B1A9),
.INIT_07(256'h1FFD25F782D9E31A88996140763BC12E30CDF99674B5B8795E793E8B46B826D8),
.INIT_08(256'h5939E2B2C74267408B274FD32B87F1FFAFCFEA18FBFBFBFBAE2BEEF9FBFBFBFB),
.INIT_09(256'hC511C52178AD2D5AA34630E54647852685FC628923DECF323A5B34C7FBFBFBFB),
.INIT_0A(256'hA3FD6E00B970CBA092002082E909E1A33A28DB5BFBFBFBFB649380E5FBFBFBFB),
.INIT_0B(256'h6B67122E007F88551A27F0FD76DD68613AD776095B40B8A32EDB8BEC7791789E),
.INIT_0C(256'h38AEAF09F049D6CDFD6555FD6F3D7383C5AD6A9014D654964F00A578FBFBFBFB),
.INIT_0D(256'h4A68667440A993D8F82907E6CE31CB96CDBCC0230F30A39C3A919EA7FBFBFBFB),
.INIT_0E(256'hD66658D8DB36400FC27C73FDCACC6BCFFDFF9909F822D70D1A3F3B8C253D4A52),
.INIT_0F(256'hE406DE0C792218E173629ABB8DC03AD5CB36026D8F4E4382A582C570BD43DD23),
.INIT_10(256'hFC232B05DAE1D90D08E918089EAD10CC689D1CF7000000004A8974A900000000),
.INIT_11(256'h1102B65446B303190B0DB443C412D3EA4E92D311341FEBC070B178A700000000),
.INIT_12(256'h48B68788E1477E37F636FECF62CC70318BC27B2C00000000245B9EFF00000000),
.INIT_13(256'h60A8F0C9881A7E03BE63361A43F2E7B94FD579FDE63716C772F5D1485CA67389),
.INIT_14(256'h4BF5612E8D59C8F3F9C7F639AECC8409FA3FD70C04BAE658FDB0782B00000000),
.INIT_15(256'hF082AA29FBE1F80DB76E173F0582B6DE7B97BF4D2BBE16837B34C89900000000),
.INIT_16(256'h0F43833E8D17EA9FAD610439331F3BF8D17BC672076A5B360123BE82598AE734),
.INIT_17(256'h2359F07B5CF25213FA2BD3F3B1820FD3E0993156A81404B8B9631FDB577EC6EF),
.INIT_18(256'h07D8D0FE211A22F6F312E3F36556EB379366E70CFBFBFBFBB1728F52FBFBFBFB),
.INIT_19(256'hEAF94DAFBD48F8E2F0F64FB83FE92811B56928EACFE4103B8B4A835CFBFBFBFB),
.INIT_1A(256'hB34D7C731ABC85CC0DCD053499378BCA703980D7FBFBFBFBDFA06504FBFBFBFB),
.INIT_1B(256'h9B530B3273E185F84598CDE1B8091C42B42E82061DCCED3C890E2AB3A75D8872),
.INIT_1C(256'hB00E9AD576A23308023C0DC255377FF201C42CF7FF411DA3064B83D0FBFBFBFB),
.INIT_1D(256'h0B7951D2001A03F64C95ECC4FE794D25806C44B6D045ED7880CF3362FBFBFBFB),
.INIT_1E(256'hF4B878C576EC1164569AFFC2C8E4C0032A803D89FC91A0CDFAD84579A2711CCF),
.INIT_1F(256'hD8A20B80A709A9E801D028084A79F4281B62CAAD53EFFF434298E420AC853D14),



	
	//===============================================================================
	
	.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),


	// The next set of INITP_xx are for the parity bits
	.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
	// The next set of INITP_xx are for "18Kb" configuration only
	.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_TDP_MACRO_inst (
	.DOA(DOA), // Output port-A data, width defined by READ_WIDTH_A parameter
	.DOB(DOB), // Output port-B data, width defined by READ_WIDTH_B parameter
	.ADDRA(ADDRA), // Input port-A address, width defined by Port A depth
	.ADDRB(ADDRB), // Input port-B address, width defined by Port B depth
	.CLKA(clk), // 1-bit input port-A clock
	.CLKB(clk), // 1-bit input port-B clock
		.DIA(8'h0), // Input port-A data, width defined by WRITE_WIDTH_A parameter
	.DIB(8'h0), // Input port-B data, width defined by WRITE_WIDTH_B parameter
	.ENA(EN), // 1-bit input port-A enable
	.ENB(EN), // 1-bit input port-B enable
	.REGCEA(EN), // 1-bit input port-A output register enable
	.REGCEB(EN), // 1-bit input port-B output register enable
	.RSTA(rst), // 1-bit input port-A reset
	.RSTB(rst), // 1-bit input port-B reset
	.WEA(1'b0), // Input port-A write enable, width defined by Port A depth
	.WEB(1'b0) // Input port-B write enable, width defined by Port B depth
);
// End of BRAM_TDP_MACRO_inst instantiation
endmodule
